module FSMParejasTotales(input rst, clk, j, output l);

	logic [2:0] contador; 
	
	

endmodule