module contador();

endmodule