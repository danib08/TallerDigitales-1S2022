module JuegoMemory();

endmodule