module memory();

endmodule