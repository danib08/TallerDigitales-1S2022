module testDeco();
	
	logic A, B, C, D, E, a, b, c, d, e, f, g;
	
	decodificador deco1(A, B, C, D, E, a, b, c, d, e, f, g);
	
	initial begin
		A = 0; B = 0; C = 0; D = 0; E = 0; #10; //P1
		A = 0; B = 0; C = 0; D = 0; E = 1; #10; //P2
		A = 0; B = 0; C = 0; D = 1; E = 0; #10; //P3
		A = 0; B = 0; C = 0; D = 1; E = 1; #10; //P4
		A = 0; B = 0; C = 1; D = 0; E = 0; #10; //P5
		A = 0; B = 0; C = 1; D = 0; E = 1; #10; //P6
		A = 0; B = 0; C = 1; D = 1; E = 0; #10; //P7
		A = 0; B = 0; C = 1; D = 1; E = 1; #10; //P8
		A = 0; B = 1; C = 0; D = 0; E = 0; #10; //P9
		A = 0; B = 1; C = 0; D = 0; E = 1; #10; //P10
		A = 0; B = 1; C = 0; D = 1; E = 0; #10; //P11
		A = 0; B = 1; C = 0; D = 1; E = 1; #10; //P12
		A = 0; B = 1; C = 1; D = 0; E = 0; #10; //P13
		A = 0; B = 1; C = 1; D = 0; E = 1; #10; //P14
		A = 0; B = 1; C = 1; D = 1; E = 0; #10; //P15
		A = 0; B = 1; C = 1; D = 1; E = 1; #10; //P16
		A = 1; B = 0; C = 0; D = 0; E = 0; #10; //P17
		A = 1; B = 0; C = 0; D = 0; E = 1; #10; //P18
		A = 1; B = 0; C = 0; D = 1; E = 0; #10; //P19
		A = 1; B = 0; C = 0; D = 1; E = 1; #10; //P20
		A = 1; B = 0; C = 1; D = 0; E = 0; #10; //P21
		A = 1; B = 0; C = 1; D = 0; E = 1; #10; //P22
		A = 1; B = 0; C = 1; D = 1; E = 0; #10; //P23
		A = 1; B = 0; C = 1; D = 1; E = 1; #10; //P24
		A = 1; B = 1; C = 0; D = 0; E = 0; #10; //P25
		A = 1; B = 1; C = 0; D = 0; E = 1; #10; //P26
		A = 1; B = 1; C = 0; D = 1; E = 0; #10; //P27
		A = 1; B = 1; C = 0; D = 1; E = 1; #10; //P28
		A = 1; B = 1; C = 1; D = 0; E = 0; #10; //P29 
		A = 1; B = 1; C = 1; D = 0; E = 1; #10; //P30
		A = 1; B = 1; C = 1; D = 1; E = 0; #10; //P31
		A = 1; B = 1; C = 1; D = 1; E = 1; #10; //P32
	end

endmodule