module vga_test ();

logic clk50MHz;
logic clk25MHz;
logic vga_hs;
logic vga_vs;
logic [7:0] vga_r;
logic [7:0] vga_g;
logic [7:0] vga_b;