module testRegisterFile();
	logic clk, we3;
	logic [3:0] ra1, ra2, ra3;
	logic [31:0] wd3, r15, rd1, rd2;
	
	

endmodule