module  Registro #(parameter n = 4) (input [n-1:0] a, b, input clk, rst, output [n-1:0] salida);
	
	


endmodule